module ALU( // @[:@3.2]
  input        clock, // @[:@4.4]
  input        reset, // @[:@5.4]
  input  [5:0] io_a, // @[:@6.4]
  input  [5:0] io_b, // @[:@6.4]
  input  [2:0] io_s, // @[:@6.4]
  output [5:0] io_y, // @[:@6.4]
  output [2:0] io_f // @[:@6.4]
);
  wire  _T_22; // @[ALU.scala 25:14:@15.4]
  wire [6:0] _T_23; // @[ALU.scala 26:26:@17.6]
  wire [5:0] _T_24; // @[ALU.scala 27:25:@19.6]
  wire [5:0] _T_25; // @[ALU.scala 27:40:@20.6]
  wire [6:0] _T_26; // @[ALU.scala 27:32:@21.6]
  wire  _T_27; // @[ALU.scala 29:20:@26.6]
  wire [6:0] _T_28; // @[ALU.scala 30:26:@28.8]
  wire [6:0] _T_29; // @[ALU.scala 30:26:@29.8]
  wire [6:0] _T_32; // @[ALU.scala 31:32:@33.8]
  wire  _T_33; // @[ALU.scala 33:20:@38.8]
  wire [5:0] _T_34; // @[ALU.scala 34:18:@40.10]
  wire  _T_35; // @[ALU.scala 35:20:@44.10]
  wire [5:0] _T_36; // @[ALU.scala 36:18:@46.12]
  wire  _T_37; // @[ALU.scala 37:20:@50.12]
  wire [5:0] _T_38; // @[ALU.scala 38:13:@52.14]
  wire  _T_39; // @[ALU.scala 39:20:@56.14]
  wire [5:0] _T_40; // @[ALU.scala 40:18:@58.16]
  wire [5:0] _GEN_0; // @[ALU.scala 39:30:@57.14]
  wire [5:0] _GEN_1; // @[ALU.scala 37:30:@51.12]
  wire [5:0] _GEN_2; // @[ALU.scala 35:29:@45.10]
  wire [5:0] _GEN_3; // @[ALU.scala 33:30:@39.8]
  wire [6:0] _GEN_4; // @[ALU.scala 29:32:@27.6]
  wire [6:0] _GEN_5; // @[ALU.scala 29:32:@27.6]
  wire [6:0] arith_result; // @[ALU.scala 25:24:@16.4]
  wire [6:0] _GEN_6; // @[ALU.scala 29:32:@27.6]
  wire [6:0] sext_result; // @[ALU.scala 25:24:@16.4]
  wire [6:0] _GEN_9; // @[ALU.scala 25:24:@16.4]
  wire  flag_zero; // @[ALU.scala 47:21:@64.4]
  wire [1:0] _T_44; // @[ALU.scala 50:32:@66.4]
  wire  _T_46; // @[ALU.scala 50:43:@67.4]
  wire  _T_49; // @[ALU.scala 50:81:@69.4]
  wire  flag_overflow; // @[ALU.scala 50:56:@70.4]
  wire  flag_carry; // @[ALU.scala 51:29:@72.4]
  wire [1:0] _T_52; // @[Cat.scala 30:58:@74.4]
  assign _T_22 = io_s == 3'h0; // @[ALU.scala 25:14:@15.4]
  assign _T_23 = io_a + io_b; // @[ALU.scala 26:26:@17.6]
  assign _T_24 = $signed(io_a); // @[ALU.scala 27:25:@19.6]
  assign _T_25 = $signed(io_b); // @[ALU.scala 27:40:@20.6]
  assign _T_26 = $signed(_T_24) + $signed(_T_25); // @[ALU.scala 27:32:@21.6]
  assign _T_27 = io_s == 3'h1; // @[ALU.scala 29:20:@26.6]
  assign _T_28 = io_a - io_b; // @[ALU.scala 30:26:@28.8]
  assign _T_29 = $unsigned(_T_28); // @[ALU.scala 30:26:@29.8]
  assign _T_32 = $signed(_T_24) - $signed(_T_25); // @[ALU.scala 31:32:@33.8]
  assign _T_33 = io_s == 3'h2; // @[ALU.scala 33:20:@38.8]
  assign _T_34 = io_a & io_b; // @[ALU.scala 34:18:@40.10]
  assign _T_35 = io_s == 3'h3; // @[ALU.scala 35:20:@44.10]
  assign _T_36 = io_a | io_b; // @[ALU.scala 36:18:@46.12]
  assign _T_37 = io_s == 3'h4; // @[ALU.scala 37:20:@50.12]
  assign _T_38 = ~ io_a; // @[ALU.scala 38:13:@52.14]
  assign _T_39 = io_s == 3'h5; // @[ALU.scala 39:20:@56.14]
  assign _T_40 = io_a ^ io_b; // @[ALU.scala 40:18:@58.16]
  assign _GEN_0 = _T_39 ? _T_40 : 6'h0; // @[ALU.scala 39:30:@57.14]
  assign _GEN_1 = _T_37 ? _T_38 : _GEN_0; // @[ALU.scala 37:30:@51.12]
  assign _GEN_2 = _T_35 ? _T_36 : _GEN_1; // @[ALU.scala 35:29:@45.10]
  assign _GEN_3 = _T_33 ? _T_34 : _GEN_2; // @[ALU.scala 33:30:@39.8]
  assign _GEN_4 = _T_27 ? _T_29 : 7'h0; // @[ALU.scala 29:32:@27.6]
  assign _GEN_5 = _T_27 ? $signed(_T_32) : $signed(7'sh0); // @[ALU.scala 29:32:@27.6]
  assign arith_result = _T_22 ? _T_23 : _GEN_4; // @[ALU.scala 25:24:@16.4]
  assign _GEN_6 = _T_27 ? arith_result : {{1'd0}, _GEN_3}; // @[ALU.scala 29:32:@27.6]
  assign sext_result = _T_22 ? $signed(_T_26) : $signed(_GEN_5); // @[ALU.scala 25:24:@16.4]
  assign _GEN_9 = _T_22 ? arith_result : _GEN_6; // @[ALU.scala 25:24:@16.4]
  assign flag_zero = io_y == 6'h0; // @[ALU.scala 47:21:@64.4]
  assign _T_44 = sext_result[6:5]; // @[ALU.scala 50:32:@66.4]
  assign _T_46 = _T_44 == 2'h1; // @[ALU.scala 50:43:@67.4]
  assign _T_49 = _T_44 == 2'h2; // @[ALU.scala 50:81:@69.4]
  assign flag_overflow = _T_46 | _T_49; // @[ALU.scala 50:56:@70.4]
  assign flag_carry = arith_result[6]; // @[ALU.scala 51:29:@72.4]
  assign _T_52 = {flag_carry,flag_overflow}; // @[Cat.scala 30:58:@74.4]
  assign io_y = _GEN_9[5:0]; // @[ALU.scala 28:10:@23.6 ALU.scala 32:10:@35.8 ALU.scala 34:10:@41.10 ALU.scala 36:10:@47.12 ALU.scala 38:10:@53.14 ALU.scala 40:10:@59.16 ALU.scala 42:10:@62.16]
  assign io_f = {_T_52,flag_zero}; // @[ALU.scala 53:8:@76.4]
endmodule

module ALU2( // @[:@3.2]
  input        clock, // @[:@4.4]
  input        reset, // @[:@5.4]
  input  [5:0] io_a, // @[:@6.4]
  input  [5:0] io_b, // @[:@6.4]
  input  [2:0] io_s, // @[:@6.4]
  output [5:0] io_y, // @[:@6.4]
  output [2:0] io_f // @[:@6.4]
);
  wire  _T_22; // @[ALU2.scala 25:14:@15.4]
  wire [6:0] _T_23; // @[ALU2.scala 26:26:@17.6]
  wire [5:0] _T_24; // @[ALU2.scala 27:25:@19.6]
  wire [5:0] _T_25; // @[ALU2.scala 27:40:@20.6]
  wire [6:0] _T_26; // @[ALU2.scala 27:32:@21.6]
  wire  _T_27; // @[ALU2.scala 29:20:@26.6]
  wire [6:0] _T_28; // @[ALU2.scala 30:26:@28.8]
  wire [6:0] _T_29; // @[ALU2.scala 30:26:@29.8]
  wire [6:0] _T_32; // @[ALU2.scala 31:32:@33.8]
  wire  _T_33; // @[ALU2.scala 33:20:@38.8]
  wire [5:0] _T_34; // @[ALU2.scala 34:18:@40.10]
  wire  _T_35; // @[ALU2.scala 35:20:@44.10]
  wire [5:0] _T_36; // @[ALU2.scala 36:18:@46.12]
  wire  _T_37; // @[ALU2.scala 37:20:@50.12]
  wire [5:0] _T_38; // @[ALU2.scala 38:13:@52.14]
  wire  _T_39; // @[ALU2.scala 39:20:@56.14]
  wire [5:0] _T_40; // @[ALU2.scala 40:18:@58.16]
  wire  _T_41; // @[ALU2.scala 41:20:@62.16]
  wire [68:0] _GEN_12; // @[ALU2.scala 42:18:@64.18]
  wire [68:0] _T_42; // @[ALU2.scala 42:18:@64.18]
  wire  _T_43; // @[ALU2.scala 43:20:@68.18]
  wire [5:0] _T_44; // @[ALU2.scala 44:18:@70.20]
  wire [5:0] _GEN_0; // @[ALU2.scala 43:29:@69.18]
  wire [68:0] _GEN_1; // @[ALU2.scala 41:29:@63.16]
  wire [68:0] _GEN_2; // @[ALU2.scala 39:30:@57.14]
  wire [68:0] _GEN_3; // @[ALU2.scala 37:30:@51.12]
  wire [68:0] _GEN_4; // @[ALU2.scala 35:29:@45.10]
  wire [68:0] _GEN_5; // @[ALU2.scala 33:30:@39.8]
  wire [6:0] _GEN_6; // @[ALU2.scala 29:32:@27.6]
  wire [6:0] _GEN_7; // @[ALU2.scala 29:32:@27.6]
  wire [6:0] arith_result; // @[ALU2.scala 25:24:@16.4]
  wire [68:0] _GEN_8; // @[ALU2.scala 29:32:@27.6]
  wire [6:0] sext_result; // @[ALU2.scala 25:24:@16.4]
  wire [68:0] _GEN_11; // @[ALU2.scala 25:24:@16.4]
  wire  flag_zero; // @[ALU2.scala 49:21:@76.4]
  wire [1:0] _T_48; // @[ALU2.scala 50:32:@78.4]
  wire  _T_50; // @[ALU2.scala 50:43:@79.4]
  wire  _T_53; // @[ALU2.scala 50:81:@81.4]
  wire  flag_overflow; // @[ALU2.scala 50:56:@82.4]
  wire  flag_carry; // @[ALU2.scala 51:29:@84.4]
  wire [1:0] _T_56; // @[Cat.scala 30:58:@86.4]
  assign _T_22 = io_s == 3'h0; // @[ALU2.scala 25:14:@15.4]
  assign _T_23 = io_a + io_b; // @[ALU2.scala 26:26:@17.6]
  assign _T_24 = $signed(io_a); // @[ALU2.scala 27:25:@19.6]
  assign _T_25 = $signed(io_b); // @[ALU2.scala 27:40:@20.6]
  assign _T_26 = $signed(_T_24) + $signed(_T_25); // @[ALU2.scala 27:32:@21.6]
  assign _T_27 = io_s == 3'h1; // @[ALU2.scala 29:20:@26.6]
  assign _T_28 = io_a - io_b; // @[ALU2.scala 30:26:@28.8]
  assign _T_29 = $unsigned(_T_28); // @[ALU2.scala 30:26:@29.8]
  assign _T_32 = $signed(_T_24) - $signed(_T_25); // @[ALU2.scala 31:32:@33.8]
  assign _T_33 = io_s == 3'h2; // @[ALU2.scala 33:20:@38.8]
  assign _T_34 = io_a & io_b; // @[ALU2.scala 34:18:@40.10]
  assign _T_35 = io_s == 3'h3; // @[ALU2.scala 35:20:@44.10]
  assign _T_36 = io_a | io_b; // @[ALU2.scala 36:18:@46.12]
  assign _T_37 = io_s == 3'h4; // @[ALU2.scala 37:20:@50.12]
  assign _T_38 = ~ io_a; // @[ALU2.scala 38:13:@52.14]
  assign _T_39 = io_s == 3'h5; // @[ALU2.scala 39:20:@56.14]
  assign _T_40 = io_a ^ io_b; // @[ALU2.scala 40:18:@58.16]
  assign _T_41 = io_s == 3'h6; // @[ALU2.scala 41:20:@62.16]
  assign _GEN_12 = {{63'd0}, io_a}; // @[ALU2.scala 42:18:@64.18]
  assign _T_42 = _GEN_12 << io_b; // @[ALU2.scala 42:18:@64.18]
  assign _T_43 = io_s == 3'h7; // @[ALU2.scala 43:20:@68.18]
  assign _T_44 = io_a >> io_b; // @[ALU2.scala 44:18:@70.20]
  assign _GEN_0 = _T_43 ? _T_44 : 6'h0; // @[ALU2.scala 43:29:@69.18]
  assign _GEN_1 = _T_41 ? _T_42 : {{63'd0}, _GEN_0}; // @[ALU2.scala 41:29:@63.16]
  assign _GEN_2 = _T_39 ? {{63'd0}, _T_40} : _GEN_1; // @[ALU2.scala 39:30:@57.14]
  assign _GEN_3 = _T_37 ? {{63'd0}, _T_38} : _GEN_2; // @[ALU2.scala 37:30:@51.12]
  assign _GEN_4 = _T_35 ? {{63'd0}, _T_36} : _GEN_3; // @[ALU2.scala 35:29:@45.10]
  assign _GEN_5 = _T_33 ? {{63'd0}, _T_34} : _GEN_4; // @[ALU2.scala 33:30:@39.8]
  assign _GEN_6 = _T_27 ? _T_29 : 7'h0; // @[ALU2.scala 29:32:@27.6]
  assign _GEN_7 = _T_27 ? $signed(_T_32) : $signed(7'sh0); // @[ALU2.scala 29:32:@27.6]
  assign arith_result = _T_22 ? _T_23 : _GEN_6; // @[ALU2.scala 25:24:@16.4]
  assign _GEN_8 = _T_27 ? {{62'd0}, arith_result} : _GEN_5; // @[ALU2.scala 29:32:@27.6]
  assign sext_result = _T_22 ? $signed(_T_26) : $signed(_GEN_7); // @[ALU2.scala 25:24:@16.4]
  assign _GEN_11 = _T_22 ? {{62'd0}, arith_result} : _GEN_8; // @[ALU2.scala 25:24:@16.4]
  assign flag_zero = io_y == 6'h0; // @[ALU2.scala 49:21:@76.4]
  assign _T_48 = sext_result[6:5]; // @[ALU2.scala 50:32:@78.4]
  assign _T_50 = _T_48 == 2'h1; // @[ALU2.scala 50:43:@79.4]
  assign _T_53 = _T_48 == 2'h2; // @[ALU2.scala 50:81:@81.4]
  assign flag_overflow = _T_50 | _T_53; // @[ALU2.scala 50:56:@82.4]
  assign flag_carry = arith_result[6]; // @[ALU2.scala 51:29:@84.4]
  assign _T_56 = {flag_carry,flag_overflow}; // @[Cat.scala 30:58:@86.4]
  assign io_y = _GEN_11[5:0]; // @[ALU2.scala 28:10:@23.6 ALU2.scala 32:10:@35.8 ALU2.scala 34:10:@41.10 ALU2.scala 36:10:@47.12 ALU2.scala 38:10:@53.14 ALU2.scala 40:10:@59.16 ALU2.scala 42:10:@65.18 ALU2.scala 44:10:@71.20 ALU2.scala 46:10:@74.20]
  assign io_f = {_T_56,flag_zero}; // @[ALU2.scala 53:8:@88.4]
endmodule

module ALU( // @[:@3.2]
  input  [5:0] io_a, // @[:@6.4]
  input  [5:0] io_b, // @[:@6.4]
  output [5:0] io_y, // @[:@6.4]
  output [2:0] io_f // @[:@6.4]
);
  wire [5:0] _T_24; // @[ALU.scala 27:25:@19.6]
  wire [5:0] _T_25; // @[ALU.scala 27:40:@20.6]
  wire [6:0] _T_28; // @[ALU.scala 30:26:@28.8]
  wire [6:0] arith_result; // @[ALU.scala 30:26:@29.8]
  wire [6:0] sext_result; // @[ALU.scala 31:32:@33.8]
  wire  flag_zero; // @[ALU.scala 47:21:@64.4]
  wire [1:0] _T_44; // @[ALU.scala 50:32:@66.4]
  wire  _T_46; // @[ALU.scala 50:43:@67.4]
  wire  _T_49; // @[ALU.scala 50:81:@69.4]
  wire  flag_overflow; // @[ALU.scala 50:56:@70.4]
  wire  flag_carry; // @[ALU.scala 51:29:@72.4]
  wire [1:0] _T_52; // @[Cat.scala 30:58:@74.4]
  assign _T_24 = $signed(io_a); // @[ALU.scala 27:25:@19.6]
  assign _T_25 = $signed(io_b); // @[ALU.scala 27:40:@20.6]
  assign _T_28 = io_a - io_b; // @[ALU.scala 30:26:@28.8]
  assign arith_result = $unsigned(_T_28); // @[ALU.scala 30:26:@29.8]
  assign sext_result = $signed(_T_24) - $signed(_T_25); // @[ALU.scala 31:32:@33.8]
  assign flag_zero = io_y == 6'h0; // @[ALU.scala 47:21:@64.4]
  assign _T_44 = sext_result[6:5]; // @[ALU.scala 50:32:@66.4]
  assign _T_46 = _T_44 == 2'h1; // @[ALU.scala 50:43:@67.4]
  assign _T_49 = _T_44 == 2'h2; // @[ALU.scala 50:81:@69.4]
  assign flag_overflow = _T_46 | _T_49; // @[ALU.scala 50:56:@70.4]
  assign flag_carry = arith_result[6]; // @[ALU.scala 51:29:@72.4]
  assign _T_52 = {flag_carry,flag_overflow}; // @[Cat.scala 30:58:@74.4]
  assign io_y = arith_result[5:0]; // @[ALU.scala 28:10:@23.6 ALU.scala 32:10:@35.8 ALU.scala 34:10:@41.10 ALU.scala 36:10:@47.12 ALU.scala 38:10:@53.14 ALU.scala 40:10:@59.16 ALU.scala 42:10:@62.16]
  assign io_f = {_T_52,flag_zero}; // @[ALU.scala 53:8:@76.4]
endmodule
module Compare( // @[:@78.2]
  input        clock, // @[:@79.4]
  input        reset, // @[:@80.4]
  input  [5:0] io_x, // @[:@81.4]
  input  [5:0] io_y, // @[:@81.4]
  output       io_ug, // @[:@81.4]
  output       io_ul, // @[:@81.4]
  output       io_eq, // @[:@81.4]
  output       io_sg, // @[:@81.4]
  output       io_sl // @[:@81.4]
);
  wire [5:0] alu_io_a; // @[Compare.scala 20:19:@83.4]
  wire [5:0] alu_io_b; // @[Compare.scala 20:19:@83.4]
  wire [5:0] alu_io_y; // @[Compare.scala 20:19:@83.4]
  wire [2:0] alu_io_f; // @[Compare.scala 20:19:@83.4]
  wire  _T_21; // @[Compare.scala 25:12:@91.4]
  wire  _T_22; // @[Compare.scala 25:30:@92.4]
  wire  _T_23; // @[Compare.scala 25:21:@93.4]
  wire  _T_29; // @[Compare.scala 27:31:@101.4]
  wire  _T_30; // @[Compare.scala 27:22:@102.4]
  wire  _T_31; // @[Compare.scala 27:49:@103.4]
  wire  _T_32; // @[Compare.scala 27:39:@104.4]
  wire  _T_37; // @[Compare.scala 28:38:@110.4]
  ALU alu ( // @[Compare.scala 20:19:@83.4]
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_y(alu_io_y),
    .io_f(alu_io_f)
  );
  assign _T_21 = ~ io_eq; // @[Compare.scala 25:12:@91.4]
  assign _T_22 = alu_io_f[2]; // @[Compare.scala 25:30:@92.4]
  assign _T_23 = ~ _T_22; // @[Compare.scala 25:21:@93.4]
  assign _T_29 = alu_io_y[5]; // @[Compare.scala 27:31:@101.4]
  assign _T_30 = ~ _T_29; // @[Compare.scala 27:22:@102.4]
  assign _T_31 = alu_io_f[1]; // @[Compare.scala 27:49:@103.4]
  assign _T_32 = _T_30 ^ _T_31; // @[Compare.scala 27:39:@104.4]
  assign _T_37 = _T_29 ^ _T_31; // @[Compare.scala 28:38:@110.4]
  assign io_ug = _T_21 & _T_23; // @[Compare.scala 25:9:@95.4]
  assign io_ul = _T_21 & _T_22; // @[Compare.scala 26:9:@99.4]
  assign io_eq = alu_io_f[0]; // @[Compare.scala 24:9:@90.4]
  assign io_sg = _T_21 & _T_32; // @[Compare.scala 27:9:@106.4]
  assign io_sl = _T_21 & _T_37; // @[Compare.scala 28:9:@112.4]
  assign alu_io_a = io_x; // @[Compare.scala 21:12:@86.4]
  assign alu_io_b = io_y; // @[Compare.scala 22:12:@87.4]
endmodule
